module onehot(din,dout);
/*
input [4:0] din;
output [4:0] dout;

reg [3:0] dout;

always @(din)

begin 
case(din)
5'b1XXXX: dout[4] <= 1;
5'b01XXX: dout[3] <= 1;
5'b001XX: dout[2] <= 1;
5'b0001x: dout[1] <= 1;
5'b00001: dout[0] <= 1;
endcase 
end 
*/
input [31:0] din;
output [31:0] dout;

reg [31:0] dout;
always @(din)
begin
case(din)
32'b1XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: dout[31] <=1;
32'b01XXXXXXXXXXXXXXXXXXXXXXXXXXXXXX: dout[30] <=1;
32'b001XXXXXXXXXXXXXXXXXXXXXXXXXXXXX: dout[29] <=1;
32'b0001XXXXXXXXXXXXXXXXXXXXXXXXXXXX: dout[28] <=1;
32'b00001XXXXXXXXXXXXXXXXXXXXXXXXXXX: dout[27] <=1;
32'b000001XXXXXXXXXXXXXXXXXXXXXXXXXX: dout[26] <=1;
32'b0000001XXXXXXXXXXXXXXXXXXXXXXXXX: dout[25] <=1;
32'b00000001XXXXXXXXXXXXXXXXXXXXXXXX: dout[24] <=1;
32'b000000001XXXXXXXXXXXXXXXXXXXXXXX: dout[23] <=1;
32'b0000000001XXXXXXXXXXXXXXXXXXXXXX: dout[22] <=1;
32'b00000000001XXXXXXXXXXXXXXXXXXXXX: dout[21] <=1;
32'b000000000001XXXXXXXXXXXXXXXXXXXX: dout[20] <=1;
32'b0000000000001XXXXXXXXXXXXXXXXXXX: dout[19] <=1;
32'b00000000000001XXXXXXXXXXXXXXXXXX: dout[18] <=1;
32'b000000000000001XXXXXXXXXXXXXXXXX: dout[17] <=1;
32'b0000000000000001XXXXXXXXXXXXXXXX: dout[16] <=1;
32'b00000000000000001XXXXXXXXXXXXXXX: dout[15] <=1;
32'b000000000000000001XXXXXXXXXXXXXX: dout[14] <=1;
32'b0000000000000000001XXXXXXXXXXXXX: dout[13] <=1;
32'b00000000000000000001XXXXXXXXXXXX: dout[12] <=1;
32'b000000000000000000001XXXXXXXXXXX: dout[11] <=1;
32'b0000000000000000000001XXXXXXXXXX: dout[10] <=1;
32'b00000000000000000000001XXXXXXXXX: dout[9] <=1;
32'b000000000000000000000001XXXXXXXX: dout[8] <=1;
32'b0000000000000000000000001XXXXXXX: dout[7] <=1;
32'b00000000000000000000000001XXXXXX: dout[6] <=1;
32'b000000000000000000000000001XXXXX: dout[5] <=1;
32'b0000000000000000000000000001XXXX: dout[4] <=1;
32'b00000000000000000000000000001XXX: dout[3] <=1;
32'b000000000000000000000000000001XX: dout[2] <=1;
32'b0000000000000000000000000000001X: dout[1] <=1;
32'b00000000000000000000000000000001: dout[0] <=1;
//32'b00000000000000000000000000000000: dout[32] <=1;

endcase
end
endmodule